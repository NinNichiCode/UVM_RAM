interface ram_if(input clk);
   logic wr;
   logic [7:0] din;
   logic [3:0] addr;
   logic [7:0] dout;

 endinterface
